<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-65.3816,-102.009,57.1566,-162.578</PageViewport>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>-24,-115.5</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-116</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>7.5,-115.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>-19,5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>-8,5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>2.5,5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>10 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>13.5,5</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>-29.5,7</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>BB_CLOCK</type>
<position>-28.5,1.5</position>
<output>
<ID>CLK</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>-13,12.5</position>
<input>
<ID>N_in2</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>-3,12.5</position>
<input>
<ID>N_in2</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>8,12.5</position>
<input>
<ID>N_in2</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>21.5,12</position>
<input>
<ID>N_in2</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-7,15.5</position>
<gparam>LABEL_TEXT 4 Bit SISO Shift Right</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-9.5,-3</position>
<gparam>LABEL_TEXT 4 Bit PISO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>-21,-30</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_DFF_LOW</type>
<position>-10.5,-30</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>47</ID>
<type>AE_DFF_LOW</type>
<position>1.5,-30</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>25 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>11,-29.5</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>50</ID>
<type>BB_CLOCK</type>
<position>-31.5,-36.5</position>
<output>
<ID>CLK</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>-18.5,-18</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>-12.5,-18</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>2.5,-18</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>9,-18</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_OR2</type>
<position>-15.5,-25</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_OR2</type>
<position>6,-24.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>-7,-18</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>-2.5,-18</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR2</type>
<position>-5,-24.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>-37.5,-9</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_INVERTER</type>
<position>-29,-9</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>-14,-6</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>-3.5,-6</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>7.5,-6</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>-33.5,-28</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>-15.5,-33</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>-4.5,-34.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>5.5,-34</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>18,-34</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>-19,-17.5</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-12.5,-17.5</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-2.5,-17.5</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>2.5,-17.5</position>
<gparam>LABEL_TEXT G5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>9,-17.5</position>
<gparam>LABEL_TEXT G6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-6.5,-17.5</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-11.5,-5.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>0,-5.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>11,-5.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>-42,-8.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-10,-45.5</position>
<gparam>LABEL_TEXT Bidirectional Shift Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AE_DFF_LOW</type>
<position>-32.5,-82</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_DFF_LOW</type>
<position>-14,-82</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_DFF_LOW</type>
<position>3.5,-82</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_DFF_LOW</type>
<position>19.5,-82</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>BB_CLOCK</type>
<position>-48.5,-85.5</position>
<output>
<ID>CLK</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND2</type>
<position>-26,-68</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>-20,-68</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_OR2</type>
<position>-23,-75</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>-26.5,-67.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>-20,-67.5</position>
<gparam>LABEL_TEXT 6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>-8,-68.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>-2,-68.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_OR2</type>
<position>-5,-75.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>-8.5,-68</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>-2,-68</position>
<gparam>LABEL_TEXT 7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_AND2</type>
<position>9,-68</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>15,-68</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_OR2</type>
<position>12,-75</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>8.5,-67.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>15,-67.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>-45,-68</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>-39,-68</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>-42,-75</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>-45.5,-67.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>-39,-67.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_TOGGLE</type>
<position>-59,-58</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_INVERTER</type>
<position>-48.5,-58</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>-60,-65.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>28.5,-64.5</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>32.5,-80</position>
<gparam>LABEL_TEXT Right O/P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>32.5,-66.5</position>
<gparam>LABEL_TEXT I/P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>-26,-81</position>
<gparam>LABEL_TEXT Left O/P</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>GA_LED</type>
<position>-23,-84.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>GA_LED</type>
<position>-4.5,-83</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>13,-84.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>29,-85</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>-15.5,-100.5</position>
<gparam>LABEL_TEXT Universal Shift Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>-61,-68.5</position>
<gparam>LABEL_TEXT I/P</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>-59.5,-52.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AE_DFF_LOW</type>
<position>-34.5,-134.5</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_DFF_LOW</type>
<position>-19,-134.5</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>156</ID>
<type>AE_DFF_LOW</type>
<position>-3,-134.5</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_DFF_LOW</type>
<position>12.5,-134.5</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_MUX_4x1</type>
<position>-35,-118.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_3</ID>71 </input>
<output>
<ID>OUT</ID>59 </output>
<input>
<ID>SEL_0</ID>64 </input>
<input>
<ID>SEL_1</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_MUX_4x1</type>
<position>-19,-118.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_3</ID>72 </input>
<output>
<ID>OUT</ID>60 </output>
<input>
<ID>SEL_0</ID>64 </input>
<input>
<ID>SEL_1</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_MUX_4x1</type>
<position>-2.5,-119</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_3</ID>73 </input>
<output>
<ID>OUT</ID>61 </output>
<input>
<ID>SEL_0</ID>64 </input>
<input>
<ID>SEL_1</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_MUX_4x1</type>
<position>12.5,-118.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>66 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>62 </output>
<input>
<ID>SEL_0</ID>64 </input>
<input>
<ID>SEL_1</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>-47,-106</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>-47,-110.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>-40,-115.5</position>
<gparam>LABEL_TEXT P1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>-24.5,-115</position>
<gparam>LABEL_TEXT P2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>-8,-115.5</position>
<gparam>LABEL_TEXT P3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>7.5,-115</position>
<gparam>LABEL_TEXT P4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>-52,-105.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>-52,-110.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>-30,-116.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>BB_CLOCK</type>
<position>-53,-141.5</position>
<output>
<ID>CLK</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_TOGGLE</type>
<position>-40,-119.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_TOGGLE</type>
<position>7.5,-121.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>27.5,-132.5</position>
<gparam>LABEL_TEXT O/P Serial SR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-40,-117</position>
<gparam>LABEL_TEXT NC</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>-24.5,-117</position>
<gparam>LABEL_TEXT NC</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-7.5,-117.5</position>
<gparam>LABEL_TEXT NC</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>7.5,-117.5</position>
<gparam>LABEL_TEXT NC</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>-44,-119</position>
<gparam>LABEL_TEXT SR I/P</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>8,-123.5</position>
<gparam>LABEL_TEXT SL I/P</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>-40,-115.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-22,-1,10.5,-1</points>
<intersection>-22 4</intersection>
<intersection>-11 3</intersection>
<intersection>-0.5 6</intersection>
<intersection>10.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11,-1,-11,4</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>-1 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-22,-1,-22,4</points>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<intersection>-1 1</intersection>
<intersection>1.5 9</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-0.5,-1,-0.5,4</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>-1 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>10.5,-1,10.5,4</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-24.5,1.5,-22,1.5</points>
<connection>
<GID>31</GID>
<name>CLK</name></connection>
<intersection>-22 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,7,-0.5,7</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-3 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-3,7,-3,11.5</points>
<connection>
<GID>35</GID>
<name>N_in2</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,7,-11,7</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-13,7,-13,11.5</points>
<connection>
<GID>33</GID>
<name>N_in2</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,7,10.5,7</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>8 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,7,8,11.5</points>
<connection>
<GID>37</GID>
<name>N_in2</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,7,-22,7</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,7,21.5,11</points>
<connection>
<GID>39</GID>
<name>N_in2</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,7,21.5,7</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,-36.5,7.5,-36.5</points>
<connection>
<GID>50</GID>
<name>CLK</name></connection>
<intersection>-23.5 4</intersection>
<intersection>-13.5 3</intersection>
<intersection>-3 7</intersection>
<intersection>7.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-13.5,-36.5,-13.5,-31</points>
<connection>
<GID>46</GID>
<name>clock</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-23.5,-36.5,-23.5,-31</points>
<intersection>-36.5 1</intersection>
<intersection>-31 14</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-3,-36.5,-3,-31</points>
<intersection>-36.5 1</intersection>
<intersection>-31 18</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>7.5,-36.5,7.5,-30.5</points>
<intersection>-36.5 1</intersection>
<intersection>-30.5 19</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-24,-31,-23.5,-31</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>-23.5 4</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-3,-31,-1.5,-31</points>
<connection>
<GID>47</GID>
<name>clock</name></connection>
<intersection>-3 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>7.5,-30.5,8,-30.5</points>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<intersection>7.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15.5,-28,-13.5,-28</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-27.5,8,-27.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-22,-16.5,-21.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-18.5,-21.5,-18.5,-21</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-18.5,-21.5,-16.5,-21.5</points>
<intersection>-18.5 1</intersection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-22,-14.5,-21.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-12.5,-21.5,-12.5,-21</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-21.5,-12.5,-21.5</points>
<intersection>-14.5 0</intersection>
<intersection>-12.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-21.5,5,-21</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-21,5,-21</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-21.5,7,-21</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,-21,9,-21</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-24,-22,-15</points>
<intersection>-24 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-24,-18,-24</points>
<intersection>-22 0</intersection>
<intersection>-18 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,-15,-19.5,-15</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,-33,-18,-24</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-33 4</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-18,-33,-16.5,-33</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-21.5,-6,-21</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7,-21,-6,-21</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-21.5,-4,-21</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4,-21,-2.5,-21</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-28,-5,-27.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-28,-1.5,-28</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-24,-10,-15</points>
<intersection>-24 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-24,-7.5,-24</points>
<intersection>-10 0</intersection>
<intersection>-7.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-15,-8,-15</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-7.5,-34.5,-7.5,-24</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 4</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-7.5,-34.5,-5.5,-34.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<intersection>-7.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-23,0,-15</points>
<intersection>-23 1</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-23,3.5,-23</points>
<intersection>0 0</intersection>
<intersection>3.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>3.5,-26.5,3.5,-23</points>
<intersection>-26.5 4</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>0,-15,1.5,-15</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>3.5,-26.5,5,-26.5</points>
<intersection>3.5 2</intersection>
<intersection>5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>5,-34,5,-26.5</points>
<intersection>-34 7</intersection>
<intersection>-28 8</intersection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>4.5,-34,5,-34</points>
<connection>
<GID>77</GID>
<name>N_in0</name></connection>
<intersection>5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>4.5,-28,5,-28</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>5 5</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35.5,-9,-32,-9</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-35 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-35,-13,-35,-9</points>
<intersection>-13 3</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-35,-13,3.5,-13</points>
<intersection>-35 2</intersection>
<intersection>-17.5 4</intersection>
<intersection>-6 6</intersection>
<intersection>3.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17.5,-15,-17.5,-13</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-13 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-6,-15,-6,-13</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-13 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>3.5,-15,3.5,-13</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-13 3</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-15,-11.5,-9</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-9,10,-9</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 0</intersection>
<intersection>-1.5 3</intersection>
<intersection>10 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-15,-1.5,-9</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>10,-15,10,-9</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-15,-13.5,-11.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-14,-11.5,-14,-8</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-11.5,-13.5,-11.5</points>
<intersection>-14 1</intersection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-15,-3.5,-8</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-15,8,-11.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>7.5,-11.5,7.5,-8</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-11.5,8,-11.5</points>
<intersection>7.5 1</intersection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31.5,-28,-24,-28</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-34,15.5,-27.5</points>
<intersection>-34 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-27.5,15.5,-27.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-34,17,-34</points>
<connection>
<GID>79</GID>
<name>N_in0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35.5,-88,16.5,-88</points>
<intersection>-35.5 4</intersection>
<intersection>-17 3</intersection>
<intersection>0.5 6</intersection>
<intersection>16.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17,-88,-17,-83</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<intersection>-88 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-35.5,-88,-35.5,-83</points>
<connection>
<GID>99</GID>
<name>clock</name></connection>
<intersection>-88 1</intersection>
<intersection>-85.5 9</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>0.5,-88,0.5,-83</points>
<connection>
<GID>101</GID>
<name>clock</name></connection>
<intersection>-88 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>16.5,-88,16.5,-83</points>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-44.5,-85.5,-35.5,-85.5</points>
<connection>
<GID>103</GID>
<name>CLK</name></connection>
<intersection>-35.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-72,-24,-71.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-26,-71.5,-26,-71</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-26,-71.5,-24,-71.5</points>
<intersection>-26 1</intersection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-72,-22,-71.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-20,-71.5,-20,-71</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-22,-71.5,-20,-71.5</points>
<intersection>-22 0</intersection>
<intersection>-20 1</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-72.5,-6,-72</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>-72 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-8,-72,-8,-71.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,-72,-6,-72</points>
<intersection>-8 1</intersection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-72.5,-4,-72</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-72 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-2,-72,-2,-71.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4,-72,-2,-72</points>
<intersection>-4 0</intersection>
<intersection>-2 1</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-72,11,-71.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9,-71.5,9,-71</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,-71.5,11,-71.5</points>
<intersection>9 1</intersection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-72,13,-71.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>15,-71.5,15,-71</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13,-71.5,15,-71.5</points>
<intersection>13 0</intersection>
<intersection>15 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-72,-43,-71.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-45,-71.5,-45,-71</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-45,-71.5,-43,-71.5</points>
<intersection>-45 1</intersection>
<intersection>-43 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41,-72,-41,-71.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-39,-71.5,-39,-71</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-41,-71.5,-39,-71.5</points>
<intersection>-41 0</intersection>
<intersection>-39 1</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-80,-42,-78</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42,-80,-35.5,-80</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-42 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-80,-23,-78</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23,-80,-17,-80</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-80,-5,-78.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-80,0.5,-80</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-80,12,-78</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-80,16.5,-80</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-65,-38,-62.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,-62.5,16,-62.5</points>
<intersection>-54.5 2</intersection>
<intersection>-38 0</intersection>
<intersection>-19 5</intersection>
<intersection>-1 7</intersection>
<intersection>16 9</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-54.5,-62.5,-54.5,-58</points>
<intersection>-62.5 1</intersection>
<intersection>-58 3</intersection>
<intersection>-58 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-57,-58,-51.5,-58</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-19,-65,-19,-62.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-1,-65.5,-1,-62.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>16,-65,16,-62.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-65,-45.5,-58</points>
<intersection>-65 4</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-58,8,-58</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 0</intersection>
<intersection>-27 3</intersection>
<intersection>-9 6</intersection>
<intersection>8 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27,-65,-27,-58</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-46,-65,-45.5,-65</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-9,-65.5,-9,-58</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>8,-65,8,-58</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-65,-40,-64</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-64,-40,-64</points>
<intersection>-58 2</intersection>
<intersection>-40 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-58,-65.5,-58,-64</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-84.5,-29,-64.5</points>
<intersection>-84.5 4</intersection>
<intersection>-80 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-80,-29,-80</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,-64.5,-21,-64.5</points>
<intersection>-29 0</intersection>
<intersection>-21 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-21,-65,-21,-64.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-29,-84.5,-24,-84.5</points>
<connection>
<GID>143</GID>
<name>N_in0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-83,-10.5,-63.5</points>
<intersection>-83 6</intersection>
<intersection>-80 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-80,-10.5,-80</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,-63.5,-3,-63.5</points>
<intersection>-44 5</intersection>
<intersection>-10.5 0</intersection>
<intersection>-3 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-3,-65.5,-3,-63.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-44,-65,-44,-63.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-10.5,-83,-5.5,-83</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-84.5,6.5,-61</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 6</intersection>
<intersection>-64 2</intersection>
<intersection>-61 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-64,14,-64</points>
<intersection>6.5 0</intersection>
<intersection>14 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-65,14,-64</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25,-61,6.5,-61</points>
<intersection>-25 5</intersection>
<intersection>6.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-25,-65,-25,-61</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-61 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>6.5,-84.5,12,-84.5</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-65.5,-7,-60</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-60,22.5,-60</points>
<intersection>-7 0</intersection>
<intersection>22.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>22.5,-85,22.5,-60</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-85 3</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-85,28,-85</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<intersection>22.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-65,10,-64.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-64.5,26.5,-64.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-141.5,9.5,-141.5</points>
<connection>
<GID>178</GID>
<name>CLK</name></connection>
<intersection>-37.5 4</intersection>
<intersection>-22 3</intersection>
<intersection>-6 6</intersection>
<intersection>9.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22,-141.5,-22,-135.5</points>
<connection>
<GID>155</GID>
<name>clock</name></connection>
<intersection>-141.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-37.5,-141.5,-37.5,-135.5</points>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<intersection>-141.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-6,-141.5,-6,-135.5</points>
<connection>
<GID>156</GID>
<name>clock</name></connection>
<intersection>-141.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>9.5,-141.5,9.5,-135.5</points>
<connection>
<GID>157</GID>
<name>clock</name></connection>
<intersection>-141.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-127.5,-32,-118.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>-127.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37.5,-127.5,-32,-127.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-37.5,-132.5,-37.5,-127.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-127.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-129,-16,-118.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-129,-16,-129</points>
<intersection>-22 2</intersection>
<intersection>-16 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-22,-132.5,-22,-129</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-129 1</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-128.5,1,-119</points>
<intersection>-128.5 1</intersection>
<intersection>-119 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-128.5,1,-128.5</points>
<intersection>-6 3</intersection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0.5,-119,1,-119</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>1 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-132.5,-6,-128.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-128.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-128.5,15.5,-118.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-128.5,15.5,-128.5</points>
<intersection>9.5 2</intersection>
<intersection>15.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9.5,-132.5,9.5,-128.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-128.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-113.5,-35,-110.5</points>
<connection>
<GID>161</GID>
<name>SEL_1</name></connection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-110.5,12.5,-110.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>-35 0</intersection>
<intersection>-19 6</intersection>
<intersection>-2.5 3</intersection>
<intersection>12.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2.5,-114,-2.5,-110.5</points>
<connection>
<GID>163</GID>
<name>SEL_1</name></connection>
<intersection>-110.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>12.5,-113.5,12.5,-110.5</points>
<connection>
<GID>164</GID>
<name>SEL_1</name></connection>
<intersection>-110.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-19,-113.5,-19,-110.5</points>
<connection>
<GID>162</GID>
<name>SEL_1</name></connection>
<intersection>-110.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-113.5,-34,-106</points>
<connection>
<GID>161</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-106,13.5,-106</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>-34 0</intersection>
<intersection>-18 6</intersection>
<intersection>-1.5 3</intersection>
<intersection>13.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-114,-1.5,-106</points>
<connection>
<GID>163</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>13.5,-113.5,13.5,-106</points>
<connection>
<GID>164</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-18,-113.5,-18,-106</points>
<connection>
<GID>162</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-126,-40,-121.5</points>
<intersection>-126 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-126,-14.5,-126</points>
<intersection>-40 0</intersection>
<intersection>-14.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-40,-121.5,-38,-121.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-132.5,-14.5,-120</points>
<intersection>-132.5 4</intersection>
<intersection>-126 1</intersection>
<intersection>-120 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-16,-132.5,-14.5,-132.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-14.5,-120,-5.5,-120</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>-14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-132.5,2,-119.5</points>
<intersection>-132.5 1</intersection>
<intersection>-123.5 2</intersection>
<intersection>-119.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-132.5,2,-132.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,-123.5,2,-123.5</points>
<intersection>-22 3</intersection>
<intersection>2 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22,-123.5,-22,-121.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>2,-119.5,9.5,-119.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-126.5,-5.5,-122</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,-126.5,17,-126.5</points>
<intersection>-5.5 0</intersection>
<intersection>17 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>17,-132.5,17,-126.5</points>
<intersection>-132.5 3</intersection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>15.5,-132.5,17,-132.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>17 2</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-132.5,-26.5,-119.5</points>
<intersection>-132.5 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31.5,-132.5,-26.5,-132.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-119.5,-22,-119.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-119.5,-38,-119.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-121.5,9.5,-121.5</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-115.5,-38,-115.5</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-115.5,-22,-115.5</points>
<connection>
<GID>162</GID>
<name>IN_3</name></connection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-115.5,-22,-115.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-116,-5.5,-116</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>163</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-115.5,9.5,-115.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<connection>
<GID>164</GID>
<name>IN_3</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>